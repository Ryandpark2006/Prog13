// module ALU(
//     input wire [4:0] opcode,
//     input wire [63:0] operand1,
//     input wire [63:0] operand2,
//     input wire [63:0] operand3,
//     input wire [63:0] signExtendedLiteral,
//     input wire [63:0] pc,
//     input wire [63:0] stackPointer,
//     input wire [63:0] memoryReadVal,
//     output reg [63:0] result,
//     output reg [63:0] readWriteAddress,
//     output reg [63:0] updated_next,
//     output reg changing_pc,
//     output reg writeEnable,
//     output reg mem_write_enable,
//     output reg halt
// );
//     always @(*) begin
//         // Default values (same as reference)
//         result            = 64'd0;
//         readWriteAddress  = 64'd0;
//         updated_next      = pc + 64'd4;
//         writeEnable       = 1'b1;
//         mem_write_enable  = 1'b0;
//         changing_pc       = 1'b0;
//         halt              = 1'b0;

//         case (opcode)
//             5'h00: result = operand1 & operand2;                         // and
//             5'h01: result = operand1 | operand2;                         // or
//             5'h02: result = operand1 ^ operand2;                         // xor
//             5'h03: result = ~operand1;                                   // not
//             5'h04: result = operand1 >> operand2[5:0];                   // shftr
//             5'h05: result = operand3 >> signExtendedLiteral;            // shftri
//             5'h06: result = operand1 << operand2[5:0];                   // shftl
//             5'h07: result = operand3 << signExtendedLiteral;            // shftli

//             5'h08: begin                                                 // br rd
//                 changing_pc  = 1;
//                 writeEnable  = 0;
//                 updated_next = operand3;
//             end
//             5'h09: begin                                                 // brr rd
//                 changing_pc  = 1;
//                 writeEnable  = 0;
//                 updated_next = pc + operand3;
//             end
//             5'h0a: begin                                                 // brr L
//                 changing_pc  = 1;
//                 writeEnable  = 0;
//                 updated_next = pc + signExtendedLiteral;
//             end
//             5'h0b: begin                                                 // brnz rd, rs
//                 writeEnable = 0;
//                 if (operand1 != 0) begin
//                     updated_next = operand3;
//                     changing_pc = 1;
//                 end
//             end
//             5'h0c: begin                                                 // call rd, rs, rt
//                 writeEnable       = 0;
//                 mem_write_enable  = 1;
//                 changing_pc       = 1;
//                 updated_next      = operand3;
//                 readWriteAddress  = stackPointer - 64'd8;
//                 result            = pc + 64'd4;
//             end
//             5'h0d: begin                                                 // return
//                 writeEnable       = 0;
//                 changing_pc       = 1;
//                 readWriteAddress  = stackPointer - 64'd8;
//                 updated_next      = memoryReadVal;
//             end
//             5'h0e: begin                                                 // brgt rd, rs, rt
//                 writeEnable = 0;
//                 if ($signed(operand1) > $signed(operand2)) begin
//                     updated_next = operand3;
//                     changing_pc = 1;
//                 end
//             end
//             5'h0f: begin                                                 // priv
//                 writeEnable = 0;
//                 if (signExtendedLiteral[3:0] == 4'h0) begin
//                     halt = 1;
//                 end
//             end
//             5'h10: begin                                                 // mov rd, (rs)(L)
//                 readWriteAddress = operand1 + signExtendedLiteral;
//                 result = memoryReadVal;
//             end
//             5'h11: result = operand1;                                    // mov rd, rs
//             5'h12: result = {operand3[63:12], signExtendedLiteral[11:0]};// mov rd, L
//             5'h13: begin                                                 // mov (rd)(L), rs
//                 writeEnable = 0;
//                 mem_write_enable = 1;
//                 readWriteAddress = operand3 + signExtendedLiteral;
//                 result = operand1;
//             end
//             5'h14: result = $realtobits($bitstoreal(operand1) + $bitstoreal(operand2)); // addf
//             5'h15: result = $realtobits($bitstoreal(operand1) - $bitstoreal(operand2)); // subf
//             5'h16: result = $realtobits($bitstoreal(operand1) * $bitstoreal(operand2)); // mulf
//             5'h17: result = $realtobits($bitstoreal(operand1) / $bitstoreal(operand2)); // divf

//             5'h18: result = operand1 + operand2;                         // add
//             5'h19: result = operand3 + signExtendedLiteral;             // addi
//             5'h1a: result = operand1 - operand2;                         // sub
//             5'h1b: result = operand3 - signExtendedLiteral;             // subi
//             5'h1c: result = operand1 * operand2;                         // mul
//             5'h1d: result = (operand2 == 0) ? 64'd0 : operand1 / operand2; // div

//             default: begin
//                 writeEnable = 0;
//                 mem_write_enable = 0;
//                 changing_pc = 0;
//             end
//         endcase
//     end
// endmodule




// module FPU(
//     input wire [63:0] operand1,
//     input wire [63:0] operand2,
//     input wire [4:0] opcode,
//     output reg [63:0] result,
//     output reg writeEnable
// );
//     always @(*) begin
//         case (opcode)
//             5'b10100: result = $realtobits($bitstoreal(operand1) + $bitstoreal(operand2));
//             5'b10101: result = $realtobits($bitstoreal(operand1) - $bitstoreal(operand2));
//             5'b10110: result = $realtobits($bitstoreal(operand1) * $bitstoreal(operand2));
//             5'b10111: result = $realtobits($bitstoreal(operand1) / $bitstoreal(operand2));
//             default:  result = 64'b0;
//         endcase
//         writeEnable = 1;
//     end
// endmodule

// module instruction_decoder(
//     input  wire [31:0] instruction,
//     output wire [4:0]  controlSignal,
//     output wire [4:0]  rd,
//     output wire [4:0]  rs,
//     output wire [4:0]  rt,
//     output wire [11:0] L,
//     output wire        rtPassed
// );
//     assign controlSignal = instruction[31:27];
//     assign rd            = instruction[26:22];
//     assign rs            = instruction[21:17];
//     assign rt            = instruction[16:12];
//     assign L             = instruction[11:0];
//     assign rtPassed = !(controlSignal == 5'b11001 ||  // addi
//                     controlSignal == 5'b11011 ||  // subi
//                     controlSignal == 5'b00101 ||  // shftri
//                     controlSignal == 5'b00111 ||  // shftli
//                     controlSignal == 5'b10010 ||  // mov_L_to_reg
//                     controlSignal == 5'b01010 ||  // brr
//                     controlSignal == 5'b10011 ||  // store
//                     controlSignal == 5'b10000);   // load

//     // assign rtPassed      = (controlSignal == 5'b11001 || controlSignal == 5'b11011 ||
//     //                         controlSignal == 5'b00101 || controlSignal == 5'b00111 ||
//     //                         controlSignal == 5'b10010 || controlSignal == 5'b01010 ||
//     //                         controlSignal == 5'b10011 || controlSignal == 5'b10000)
//     //                        ? 0 : 1;
// endmodule

// module memory(
//     input  wire [63:0] pc,
//     input  wire        clk,
//     input  wire        reset,
//     input  wire        mem_write_enable,
//     input  wire [63:0] rw_val,
//     input  wire [31:0] rw_addr,
//     output wire [31:0] instruction,
//     output wire [63:0] r_out
// );
//     reg [7:0] bytes [524287:0];

//     assign instruction = {bytes[pc+3], bytes[pc+2], bytes[pc+1], bytes[pc]};
//     assign r_out       = {bytes[rw_addr+7], bytes[rw_addr+6], bytes[rw_addr+5], bytes[rw_addr+4],
//                           bytes[rw_addr+3], bytes[rw_addr+2], bytes[rw_addr+1], bytes[rw_addr]};

//     integer i;
//     always @(posedge clk or posedge reset) begin
//         if (reset) begin
//             for (i = 0; i < 524288; i = i + 1)
//                 bytes[i] <= 8'b0;
//         end else if (mem_write_enable) begin
//             bytes[rw_addr+7] <= rw_val[63:56];
//             bytes[rw_addr+6] <= rw_val[55:48];
//             bytes[rw_addr+5] <= rw_val[47:40];
//             bytes[rw_addr+4] <= rw_val[39:32];
//             bytes[rw_addr+3] <= rw_val[31:24];
//             bytes[rw_addr+2] <= rw_val[23:16];
//             bytes[rw_addr+1] <= rw_val[15:8];
//             bytes[rw_addr  ] <= rw_val[7:0];
//         end
//     end
// endmodule

// module register_file(
//     input  wire        clk,
//     input  wire        reset,
//     input  wire        write_enable,
//     input  wire [63:0] dataInput,
//     input  wire [4:0]  readAddress1,
//     input  wire [4:0]  readAddress2,
//     input  wire [4:0]  readAddress3,
//     input  wire [4:0]  writeAddress,
//     input  wire        lPassed,
//     input  wire [11:0] L,
//     output wire [63:0] value1,
//     output wire [63:0] value2,
//     output wire [63:0] rdVal,
//     output wire [63:0] r31_val
// );
//     reg [63:0] registers [31:0];

//     assign value1 = registers[readAddress1];
//     assign value2 = lPassed ? {{52{L[11]}},L} : registers[readAddress2];
//     assign rdVal  = registers[readAddress3];
//     assign r31_val= registers[31];

//     integer j;
//     always @(posedge clk) begin
//         if (reset) begin
//             for (j = 0; j < 31; j = j + 1)
//                 registers[j] <= 64'b0;
//             registers[31] <= 64'h80000;
//         end else if (write_enable) begin
//             registers[writeAddress] <= dataInput;
//         end
//     end
// endmodule

// module tinker_core(
//     input  wire        clk,
//     input  wire        reset,
//     output wire        hlt
// );
//     reg [63:0] PC;
//     reg [1:0]  stall_cnt;

//     reg [63:0] IF_ID_PC;
//     reg [31:0] IF_ID_IR;

//     wire [4:0]  IF_ctrl, IF_rd, IF_rs, IF_rt;
//     wire [11:0] IF_L;
//     wire        IF_rtPassed;

//     instruction_decoder dec(
//         .instruction  (IF_ID_IR),
//         .controlSignal(IF_ctrl),
//         .rd           (IF_rd),
//         .rs           (IF_rs),
//         .rt           (IF_rt),
//         .L            (IF_L),
//         .rtPassed     (IF_rtPassed)
//     );

//     wire load_use_hazard = (EX_MEM_ctrl == 5'b10000) && (
//         (IF_ctrl != 5'h1F && EX_MEM_rd == IF_rs) ||
//         (IF_ctrl != 5'h1F && EX_MEM_rd == IF_rt && IF_rtPassed)
//     );

//     wire flushFetch = aluChangePC;
//     wire fetchStall = load_use_hazard || (stall_cnt != 0);

//     wire [31:0] inst;
//     wire [63:0] mem_rdata;
//     memory memory (
//         .pc               (PC),
//         .clk              (clk),
//         .reset            (reset),
//         .mem_write_enable (EX_MEM_memWrite),
//         .rw_val           (EX_MEM_wrData),
//         .rw_addr          (EX_MEM_addr[31:0]),
//         .instruction      (inst),
//         .r_out            (mem_rdata)
//     );

//     wire [31:0] next_IF_ID_IR = flushFetch ? 32'd0 :
//                                 fetchStall ? IF_ID_IR :
//                                              inst;
//     wire [63:0] next_IF_ID_PC = flushFetch ? 64'd0 :
//                                 fetchStall ? IF_ID_PC :
//                                              PC;

//     reg [63:0] ID_EX_PC;
//     reg [4:0]  ID_EX_ctrl, ID_EX_rd, ID_EX_rs, ID_EX_rt;
//     reg [11:0] ID_EX_L;
//     reg        ID_EX_rtPassed;
//     reg [63:0] ID_EX_A, ID_EX_B;
//     reg [63:0] ID_EX_r31, ID_EX_rdVal;

//     reg [4:0]  EX_MEM_ctrl, EX_MEM_rd;
//     reg [63:0] EX_MEM_ALU, EX_MEM_B;
//     reg        EX_MEM_memWrite, EX_MEM_regWrite, EX_MEM_changePC;
//     reg [63:0] EX_MEM_addr, EX_MEM_wrData, EX_MEM_target;

//     reg [4:0]  MEM_WB_ctrl, MEM_WB_rd;
//     reg [63:0] MEM_WB_ALU, MEM_WB_memData;
//     reg        MEM_WB_regWrite, MEM_WB_memToReg;

//     wire [63:0] regOut1, regOut2, rdValSignal, r31Val;
//     register_file reg_file(
//         .clk         (clk),
//         .reset       (reset),
//         .write_enable(MEM_WB_regWrite),
//         .dataInput   (MEM_WB_memToReg ? MEM_WB_memData : MEM_WB_ALU),
//         .readAddress1(IF_rs),
//         .readAddress2(IF_rt),
//         .readAddress3(IF_rd),
//         .writeAddress(MEM_WB_rd),
//         .lPassed     (~IF_rtPassed),
//         .L           (IF_L),
//         .value1      (regOut1),
//         .value2      (regOut2),
//         .rdVal       (rdValSignal),
//         .r31_val     (r31Val)
//     );

//     wire forwardA_EX = EX_MEM_regWrite && (EX_MEM_rd != 0) && (EX_MEM_rd == ID_EX_rs);
//     wire forwardA_MEM = MEM_WB_regWrite && (MEM_WB_rd != 0) && (MEM_WB_rd == ID_EX_rs);
//     wire forwardB_EX = EX_MEM_regWrite && (EX_MEM_rd != 0) && (EX_MEM_rd == ID_EX_rt) && ID_EX_rtPassed;
//     wire forwardB_MEM = MEM_WB_regWrite && (MEM_WB_rd != 0) && (MEM_WB_rd == ID_EX_rt) && ID_EX_rtPassed;
//     wire forwardRD_EX = EX_MEM_regWrite && (EX_MEM_rd != 0) && (EX_MEM_rd == ID_EX_rd);
//     wire forwardRD_MEM = MEM_WB_regWrite && (MEM_WB_rd != 0) && (MEM_WB_rd == ID_EX_rd);

//     wire [63:0] forwarded_A = forwardA_EX ? EX_MEM_ALU :
//                              (forwardA_MEM ? (MEM_WB_memToReg ? MEM_WB_memData : MEM_WB_ALU) : ID_EX_A);

//     wire [63:0] forwarded_B = forwardB_EX ? EX_MEM_ALU :
//                              (forwardB_MEM ? (MEM_WB_memToReg ? MEM_WB_memData : MEM_WB_ALU) : ID_EX_B);

//     wire [63:0] forwarded_rdVal = forwardRD_EX ? EX_MEM_ALU :
//                                  (forwardRD_MEM ? (MEM_WB_memToReg ? MEM_WB_memData : MEM_WB_ALU) : ID_EX_rdVal);

//     wire [63:0] aluOp1 = (ID_EX_ctrl == 5'b11001 || ID_EX_ctrl == 5'b11011)
//                         ? forwarded_rdVal : forwarded_A;
//     wire [63:0] aluOp2 = ID_EX_rtPassed
//                         ? forwarded_B
//                         : {{52{ID_EX_L[11]}}, ID_EX_L};

//     wire [63:0] aluResult, aluAddr, aluUpdatedNext;
//     wire        aluRegWrite, aluMemWrite, aluChangePC, aluHalt;
//     ALU ALU_INST(
//         .opcode           (ID_EX_ctrl),
//         .operand1         (aluOp1),
//         .operand2         (aluOp2),
//         .operand3         (forwarded_rdVal),
//         .signExtendedLiteral({{52{ID_EX_L[11]}}, ID_EX_L}),
//         .pc               (ID_EX_PC),
//         .stackPointer     (ID_EX_r31),
//         .memoryReadVal    (mem_rdata),
//         .result           (aluResult),
//         .readWriteAddress (aluAddr),
//         .updated_next     (aluUpdatedNext),
//         .changing_pc      (aluChangePC),
//         .writeEnable      (aluRegWrite),
//         .mem_write_enable (aluMemWrite),
//         .halt             (aluHalt)
//     );

//     always @(posedge clk or posedge reset) begin
//         if (reset) begin
//             stall_cnt <= 0;
//         end else if (load_use_hazard) begin
//             stall_cnt <= 2;
//         end else if (stall_cnt != 0) begin
//             stall_cnt <= stall_cnt - 1;
//         end
//     end

//     reg halt_flag;
//     always @(posedge clk or posedge reset) begin
//         if (reset) begin
//             halt_flag <= 0;
//         end else if (aluHalt) begin
//             halt_flag <= 1;
//         end
//     end
//     assign hlt = halt_flag;

//     always @(posedge clk or posedge reset) begin
//         if (reset) begin
//             PC        <= 64'h2000;
//             IF_ID_PC  <= 0;
//             IF_ID_IR  <= 0;
//         end else begin
//             if (flushFetch)
//                 PC <= aluUpdatedNext;
//             else if (!fetchStall)
//                 PC <= PC + 4;
//             IF_ID_PC <= next_IF_ID_PC;
//             IF_ID_IR <= next_IF_ID_IR;
//         end
//     end

//     always @(posedge clk or posedge reset) begin
//         if (reset || flushFetch || fetchStall) begin
//             ID_EX_ctrl     <= 5'h1F;
//             ID_EX_rd       <= IF_rd;
//             ID_EX_rs       <= IF_rs;
//             ID_EX_rt       <= IF_rt;
//             ID_EX_L        <= IF_L;
//             ID_EX_rtPassed <= IF_rtPassed;
//             ID_EX_A        <= regOut1;
//             ID_EX_B        <= regOut2;
//             ID_EX_PC       <= IF_ID_PC;
//             ID_EX_r31      <= r31Val;
//             ID_EX_rdVal    <= rdValSignal;
//         end else begin
//             ID_EX_ctrl     <= IF_ctrl;
//             ID_EX_rd       <= IF_rd;
//             ID_EX_rs       <= IF_rs;
//             ID_EX_rt       <= IF_rt;
//             ID_EX_L        <= IF_L;
//             ID_EX_rtPassed <= IF_rtPassed;
//             ID_EX_A        <= regOut1;
//             ID_EX_B        <= regOut2;
//             ID_EX_PC       <= IF_ID_PC;
//             ID_EX_r31      <= r31Val;
//             ID_EX_rdVal    <= rdValSignal;
//         end
//     end

//     always @(posedge clk or posedge reset) begin
//         if (reset) begin
//             EX_MEM_ctrl     <= 0;
//             EX_MEM_rd       <= 0;
//             EX_MEM_ALU      <= 0;
//             EX_MEM_B        <= 0;
//             EX_MEM_memWrite <= 0;
//             EX_MEM_regWrite <= 0;
//             EX_MEM_addr     <= 0;
//             EX_MEM_wrData   <= 0;
//             EX_MEM_changePC <= 0;
//             EX_MEM_target   <= 0;
//         end else begin
//             EX_MEM_ctrl     <= ID_EX_ctrl;
//             EX_MEM_rd       <= ID_EX_rd;
//             EX_MEM_ALU      <= aluResult;
//             EX_MEM_B        <= ID_EX_B;
//             EX_MEM_memWrite <= aluMemWrite;
//             EX_MEM_regWrite <= aluRegWrite;
//             EX_MEM_addr     <= aluAddr;
//             EX_MEM_wrData   <= aluResult;
//             EX_MEM_changePC <= aluChangePC;
//             EX_MEM_target   <= aluUpdatedNext;
//         end
//     end

//     always @(posedge clk or posedge reset) begin
//         if (reset) begin
//             MEM_WB_ctrl     <= 0;
//             MEM_WB_rd       <= 0;
//             MEM_WB_ALU      <= 0;
//             MEM_WB_memData  <= 0;
//             MEM_WB_regWrite <= 0;
//             MEM_WB_memToReg <= 0;
//         end else begin
//             MEM_WB_ctrl     <= EX_MEM_ctrl;
//             MEM_WB_rd       <= EX_MEM_rd;
//             MEM_WB_ALU      <= EX_MEM_ALU;
//             MEM_WB_memData  <= mem_rdata;
//             MEM_WB_regWrite <= EX_MEM_regWrite;
//             MEM_WB_memToReg <= (EX_MEM_ctrl == 5'b10000);
//         end
//     end
// endmodule

module ALU(
    input  wire [4:0]  opcode,
    input  wire [63:0] inputDataOne,
    input  wire [63:0] inputDataTwo,
    input  wire [63:0] inputDataThree,
    input  wire [63:0] signExtendedLiteral,
    input  wire [63:0] programCounter,
    input  wire [63:0] stackPointer,
    input  wire [63:0] readMemory,
    output reg  [63:0] result,
    output reg  [63:0] readWriteAddress,
    output reg  [63:0] newProgramCounter,
    output reg         branchTaken,
    output reg         writeToRegister,
    output reg         writeToMemory,
    output reg         hlt
);
    always @(*) begin
        // ---- defaults --------------------------------------------------
        result            = 64'd0;
        readWriteAddress  = 64'd0;
        newProgramCounter = programCounter + 64'd4;
        writeToRegister   = 1'b1;
        writeToMemory     = 1'b0;
        branchTaken       = 1'b0;
        hlt               = 1'b0;
        // ---- opcode decode --------------------------------------------
        case (opcode)
            5'h00: result = inputDataOne &  inputDataTwo;                       // and
            5'h01: result = inputDataOne |  inputDataTwo;                       // or
            5'h02: result = inputDataOne ^  inputDataTwo;                       // xor
            5'h03: result = ~inputDataOne;                                      // not
            5'h04: result = inputDataOne >> inputDataTwo[5:0];                  // shftr
            5'h05: result = inputDataThree >> signExtendedLiteral;              // shftri
            5'h06: result = inputDataOne << inputDataTwo[5:0];                  // shftl
            5'h07: result = inputDataThree << signExtendedLiteral;              // shftli

            5'h08: begin                                                        // br rd
                branchTaken       = 1;
                writeToRegister   = 0;
                newProgramCounter = inputDataThree;
            end
            5'h09: begin                                                        // brr rd
                branchTaken       = 1;
                writeToRegister   = 0;
                newProgramCounter = programCounter + inputDataThree;
            end
            5'h0a: begin                                                        // brr L
                branchTaken       = 1;
                writeToRegister   = 0;
                newProgramCounter = programCounter + signExtendedLiteral;
            end
            5'h0b: begin                                                        // brnz rd,rs
                writeToRegister   = 0;
                if (inputDataOne != 64'd0) begin
                    newProgramCounter = inputDataThree;
                    branchTaken       = 1;
                end
            end
            5'h0c: begin                                                        // call rd,rs,rt
                writeToRegister   = 0;
                writeToMemory     = 1;
                branchTaken       = 1;
                newProgramCounter = inputDataThree;
                readWriteAddress  = stackPointer - 64'd8;
                result            = programCounter + 64'd4; // link
            end
            5'h0d: begin                                                        // return
                writeToRegister   = 0;
                branchTaken       = 1;
                readWriteAddress  = stackPointer - 64'd8;
                newProgramCounter = readMemory; // value popped from stack
            end
            5'h0e: begin                                                        // brgt
                writeToRegister = 0;
                if ($signed(inputDataOne) > $signed(inputDataTwo)) begin
                    newProgramCounter = inputDataThree;
                    branchTaken       = 1;
                end
            end
            5'h0f: begin                                                        // priv / halt
                writeToRegister = 0;
                if (signExtendedLiteral[3:0] == 4'h0) hlt = 1;
            end
            5'h10: begin                                                        // load  rd, (rs)(L)
                readWriteAddress  = inputDataOne + signExtendedLiteral;
                result            = readMemory;
            end
            5'h11: result = inputDataOne;                                       // mov rd,rs
            5'h12: result = {inputDataThree[63:12], signExtendedLiteral[11:0]}; // mov rd,L
            5'h13: begin                                                        // store (rd)(L),rs
                writeToRegister  = 0;
                writeToMemory    = 1;
                readWriteAddress = inputDataThree + signExtendedLiteral;
                result           = inputDataOne;
            end
            5'h14: result = $realtobits($bitstoreal(inputDataOne) + $bitstoreal(inputDataTwo)); // addf
            5'h15: result = $realtobits($bitstoreal(inputDataOne) - $bitstoreal(inputDataTwo)); // subf
            5'h16: result = $realtobits($bitstoreal(inputDataOne) * $bitstoreal(inputDataTwo)); // mulf
            5'h17: result = $realtobits($bitstoreal(inputDataOne) / $bitstoreal(inputDataTwo)); // divf

            5'h18: result = inputDataOne + inputDataTwo;                        // add
            5'h19: result = inputDataThree + signExtendedLiteral;               // addi
            5'h1a: result = inputDataOne - inputDataTwo;                        // sub
            5'h1b: result = inputDataThree - signExtendedLiteral;               // subi
            5'h1c: result = inputDataOne * inputDataTwo;                        // mul
            5'h1d: result = (inputDataTwo == 0) ? 64'd0 : (inputDataOne / inputDataTwo); // div

            default: begin
                writeToRegister = 0;
                writeToMemory   = 0;
                branchTaken     = 0;
            end
        endcase
    end
endmodule

// ===================== 2. Instruction Decoder ===============
// Interface unchanged from the original design so the register
// file keeps working the same way. We only re‑implemented the
// internals for clarity.
module instruction_decoder(
    input  wire [31:0] instruction,
    output wire [4:0]  controlSignal,
    output wire [4:0]  rd,
    output wire [4:0]  rs,
    output wire [4:0]  rt,
    output wire [11:0] L,
    output wire        rtPassed
);
    assign controlSignal = instruction[31:27];
    assign rd            = instruction[26:22];
    assign rs            = instruction[21:17];
    assign rt            = instruction[16:12];
    assign L             = instruction[11:0];

    // Immediate‑style ops do NOT forward the rt register
    assign rtPassed = !(controlSignal == 5'h19 || // addi
                         controlSignal == 5'h1b || // subi
                         controlSignal == 5'h05 || // shftri
                         controlSignal == 5'h07 || // shftli
                         controlSignal == 5'h10 || // load
                         controlSignal == 5'h0a || // brr L
                         controlSignal == 5'h13 || // store
                         controlSignal == 5'h00);  // and (literal form)
endmodule

// ===================== 3. Register File =====================
// Same external contract (so existing wrapper code keeps
// compiling) but we upgraded the internals to match reference
// behaviour (e.g. deterministic stack‑pointer initialisation).
module register_file(
    input  wire        clk,
    input  wire        reset,
    input  wire        write_enable,
    input  wire [63:0] dataInput,
    input  wire [4:0]  readAddress1,
    input  wire [4:0]  readAddress2,
    input  wire [4:0]  readAddress3,
    input  wire [4:0]  writeAddress,
    input  wire        lPassed,
    input  wire [11:0] L,
    output wire [63:0] value1,
    output wire [63:0] value2,
    output wire [63:0] rdVal,
    output wire [63:0] r31_val
);
    reg [63:0] regs [0:31];
    assign value1  = regs[readAddress1];
    assign value2  = lPassed ? {{52{L[11]}},L} : regs[readAddress2];
    assign rdVal   = regs[readAddress3];
    assign r31_val = regs[31];

    integer i;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            for (i = 0; i < 31; i = i + 1) regs[i] <= 64'd0;
            regs[31] <= 64'd524288; // stack base
        end else if (write_enable && writeAddress != 5'd0) begin
            regs[writeAddress] <= dataInput;
        end
    end
endmodule

// ===================== 4. Unified Instruction / Data Memory =
// API kept identical to the original so nothing outside this
// file needs to change.
module memory(
    input  wire        clk,
    input  wire [63:0] pc,
    input  wire        reset,
    input  wire        mem_write_enable,
    input  wire [63:0] rw_val,
    input  wire [31:0] rw_addr,
    output wire [31:0] instruction,
    output wire [63:0] r_out
);
    reg [7:0] mem [0:524287];

    assign instruction = {mem[pc+3], mem[pc+2], mem[pc+1], mem[pc  ]};
    assign r_out       = {mem[rw_addr+7], mem[rw_addr+6], mem[rw_addr+5], mem[rw_addr+4],
                          mem[rw_addr+3], mem[rw_addr+2], mem[rw_addr+1], mem[rw_addr  ]};

    integer k;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            for (k = 0; k < 524288; k = k + 1) mem[k] <= 8'd0;
        end else if (mem_write_enable) begin
            {mem[rw_addr+7], mem[rw_addr+6], mem[rw_addr+5], mem[rw_addr+4],
             mem[rw_addr+3], mem[rw_addr+2], mem[rw_addr+1], mem[rw_addr  ]} <= rw_val;
        end
    end
endmodule

// ===================== 5. Tinker Core =======================
// The pipeline has been completely rewritten. We keep the same
// observable behaviour but the control‑path is now in lock‑step
// with the course reference.
module tinker_core(
    input  wire clk,
    input  wire reset,
    output wire hlt
);
/* =============================================================
   0. Program Counter / FETCH stage ---------------------------*/
reg  [63:0] pcReg;             // current PC
wire [63:0] pcPlus4 = pcReg + 64'd4;

/* =============================================================
   1. IF / ID pipeline reg -----------------------------------*/
reg [31:0] if_id_instr;
reg [63:0] if_id_pcPlus4;

/* =============================================================
   2. ID / EX pipeline reg -----------------------------------*/
reg [4:0]  id_ex_op, id_ex_rd, id_ex_rs, id_ex_rt;
reg [63:0] id_ex_A,  id_ex_B,  id_ex_C;
reg [63:0] id_ex_seLit, id_ex_pcPlus4, id_ex_sp;
reg        id_ex_rtPassed;

/* =============================================================
   3. EX / MEM pipeline reg ----------------------------------*/
reg [4:0]  ex_mem_rd;
reg [63:0] ex_mem_result, ex_mem_addr, ex_mem_newPC;
reg        ex_mem_branch, ex_mem_wrReg, ex_mem_wrMem, ex_mem_hlt;

/* =============================================================
   4. MEM / WB pipeline reg ----------------------------------*/
reg [4:0]  mem_wb_rd;
reg [63:0] mem_wb_result;
reg        mem_wb_wrReg, mem_wb_hlt;

assign hlt = mem_wb_hlt;

/* =============================================================
   Instruction / Data memory ---------------------------------*/
wire [31:0] fetchedInstr;
wire [63:0] memReadData;

memory memory(
    .clk              (clk),
    .pc               (pcReg),
    .reset            (reset),
    .mem_write_enable (ex_mem_wrMem),
    .rw_val           (ex_mem_result), // store data
    .rw_addr          (ex_mem_addr[31:0]),
    .instruction      (fetchedInstr),
    .r_out            (memReadData)
);

/* =============================================================
   Decode -----------------------------------------------------*/
wire [4:0] op_dec, rd_dec, rs_dec, rt_dec;  wire [11:0] l_dec;  wire rtPassed_dec;

instruction_decoder DEC(
    .instruction (if_id_instr),
    .controlSignal(op_dec), .rd(rd_dec), .rs(rs_dec), .rt(rt_dec),
    .L(l_dec), .rtPassed(rtPassed_dec)
);

wire [63:0] seLiteral = {{52{l_dec[11]}}, l_dec};

/* Register file */
wire [63:0] regA, regB, regC, stackPtr;

register_file reg_file(
    .clk          (clk), .reset(reset),
    .write_enable (mem_wb_wrReg),
    .dataInput    (mem_wb_result),
    .readAddress1 (rs_dec), .readAddress2(rt_dec), .readAddress3(rd_dec),
    .writeAddress (mem_wb_rd),
    .lPassed      (~rtPassed_dec), .L(l_dec),
    .value1       (regA), .value2(regB), .rdVal(regC), .r31_val(stackPtr)
);

/* =============================================================
   5. Simple RAW hazard detector ------------------------------*/
function automatic isWriteReg(input [4:0] op);
    begin
        case (op)
            5'h08,5'h09,5'h0a,5'h0b,5'h0c,5'h0d,5'h0e,5'h0f,5'h13,5'h1F: isWriteReg = 0; // CTR‑flow, store, bubble
            default:                   isWriteReg = 1;
        endcase
    end
endfunction

wire hazard_IDEX = isWriteReg(id_ex_op) &&
                   ((id_ex_rd == rs_dec) || (id_ex_rd == rt_dec) || (id_ex_rd == rd_dec));

wire hazard_EX = ex_mem_wrReg &&
                 ((ex_mem_rd == rs_dec) || (ex_mem_rd == rt_dec) || (ex_mem_rd == rd_dec));

wire hazard_MEM = mem_wb_wrReg &&
                  ((mem_wb_rd == rs_dec) || (mem_wb_rd == rt_dec) || (mem_wb_rd == rd_dec));

wire fetchStall  = hazard_IDEX | hazard_EX | hazard_MEM;

/* =============================================================
   6. Branch flush detection ----------------------------------*/
wire alu_branchTaken;

/* =============================================================
   7. Next‑state (IF/ID) --------------------------------------*/
wire [31:0] next_if_instr   = (alu_branchTaken) ? 32'd0 : (fetchStall ? if_id_instr   : fetchedInstr);
wire [63:0] next_if_pcPlus4 = (alu_branchTaken) ? 64'd0 : (fetchStall ? if_id_pcPlus4 : pcPlus4);

/* =============================================================
   8. ALU input muxes -----------------------------------------*/
wire [63:0] aluIn1 = regA;
wire [63:0] aluIn2 = rtPassed_dec ? regB : seLiteral;
wire [63:0] aluIn3 = regC;

/* =============================================================
   9. ALU instance -------------------------------------------*/
wire [63:0] aluResult, aluAddr, aluNewPC;
wire        aluWriteReg, aluWriteMem, aluHalt;

ALU ALU_I(
    .opcode              (id_ex_op),
    .inputDataOne        (aluIn1),
    .inputDataTwo        (aluIn2),
    .inputDataThree      (aluIn3),
    .signExtendedLiteral (seLiteral),
    .programCounter      (if_id_pcPlus4 - 64'd4), // PC of current instr
    .stackPointer        (stackPtr),
    .readMemory          (memReadData),
    .result              (aluResult),
    .readWriteAddress    (aluAddr),
    .newProgramCounter   (aluNewPC),
    .branchTaken         (alu_branchTaken),
    .writeToRegister     (aluWriteReg),
    .writeToMemory       (aluWriteMem),
    .hlt                 (aluHalt)
);

/* =============================================================
   10. Sequential logic ---------------------------------------*/
localparam [4:0] BUBBLE_OP = 5'h1F;  wire bubble = fetchStall | alu_branchTaken;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        // PC & IF/ID
        pcReg           <= 64'h2000;
        if_id_instr     <= 32'd0;
        if_id_pcPlus4   <= 64'd0;
        // ID/EX
        id_ex_op        <= BUBBLE_OP;
        id_ex_rd        <= 5'd0;
        id_ex_rs        <= 5'd0;
        id_ex_rt        <= 5'd0;
        id_ex_A         <= 64'd0;
        id_ex_B         <= 64'd0;
        id_ex_C         <= 64'd0;
        id_ex_seLit     <= 64'd0;
        id_ex_pcPlus4   <= 64'd0;
        id_ex_sp        <= 64'd0;
        id_ex_rtPassed  <= 1'b0;
        // EX/MEM
        ex_mem_rd       <= 5'd0;
        ex_mem_result   <= 64'd0;
        ex_mem_addr     <= 64'd0;
        ex_mem_newPC    <= 64'd0;
        ex_mem_branch   <= 1'b0;
        ex_mem_wrReg    <= 1'b0;
        ex_mem_wrMem    <= 1'b0;
        ex_mem_hlt      <= 1'b0;
        // MEM/WB
        mem_wb_rd       <= 5'd0;
        mem_wb_result   <= 64'd0;
        mem_wb_wrReg    <= 1'b0;
        mem_wb_hlt      <= 1'b0;
    end else begin
        /* PC update */
        if (alu_branchTaken)      pcReg <= aluNewPC;
        else if (!fetchStall)     pcReg <= pcPlus4;

        /* IF/ID */
        if_id_instr   <= next_if_instr;
        if_id_pcPlus4 <= next_if_pcPlus4;

        /* ID/EX (bubble injection) */
        if (bubble) begin
            id_ex_op <= BUBBLE_OP;
        end else begin
            id_ex_op <= op_dec;
        end
        id_ex_rd       <= rd_dec;
        id_ex_rs       <= rs_dec;
        id_ex_rt       <= rt_dec;
        id_ex_A        <= regA;
        id_ex_B        <= regB;
        id_ex_C        <= regC;
        id_ex_seLit    <= seLiteral;
        id_ex_pcPlus4  <= if_id_pcPlus4;
        id_ex_sp       <= stackPtr;
        id_ex_rtPassed <= rtPassed_dec;

        /* EX/MEM */
        ex_mem_rd       <= id_ex_rd;
        ex_mem_result   <= aluResult;
        ex_mem_addr     <= aluAddr;
        ex_mem_newPC    <= aluNewPC;
        ex_mem_branch   <= alu_branchTaken;
        ex_mem_wrReg    <= aluWriteReg;
        ex_mem_wrMem    <= aluWriteMem;
        ex_mem_hlt      <= aluHalt;

        /* MEM/WB */
        mem_wb_rd     <= ex_mem_rd;
        mem_wb_result <= ex_mem_result;
        mem_wb_wrReg  <= ex_mem_wrReg;
        mem_wb_hlt    <= ex_mem_hlt;
    end
end
endmodule

// ===================== 6. Optional FPU ======================
// Retained unmodified for compatibility with any standalone
// floating‑point tests the user might have.
module FPU(
    input  wire [63:0] operand1,
    input  wire [63:0] operand2,
    input  wire [4:0]  opcode,
    output reg  [63:0] result,
    output reg         writeEnable
);
    always @(*) begin
        case (opcode)
            5'b10100: result = $realtobits($bitstoreal(operand1) + $bitstoreal(operand2));
            5'b10101: result = $realtobits($bitstoreal(operand1) - $bitstoreal(operand2));
            5'b10110: result = $realtobits($bitstoreal(operand1) * $bitstoreal(operand2));
            5'b10111: result = $realtobits($bitstoreal(operand1) / $bitstoreal(operand2));
            default:  result = 64'd0;
        endcase
        writeEnable = 1'b1;
    end
endmodule
